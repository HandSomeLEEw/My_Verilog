`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/05/08 10:19:20
// Design Name: 
// Module Name: decode_416
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module decode_416(
input [3:0] s,
output [15:0] y
    );
reg [15:0] y;

always @(s) 
begin 
	case (s)
		4'b0000:y=16'b0000_0000_0000_0001;

		4'b0001:y=16'b0000_0000_0000_0010;

		4'b0010:y=16'b0000_0000_0000_0100;

		4'b0011:y=16'b0000_0000_0000_1000;

		4'b0100:y=16'b0000_0000_0001_0000;

		4'b0101:y=16'b0000_0000_0010_0000;

		4'b0110:y=16'b0000_0000_0100_0000;

		4'b0111:y=16'b0000_0000_1000_0000;

		4'b1000:y=16'b0000_0001_0000_0000;

		4'b1001:y=16'b0000_0010_0000_0000;

		4'b1010:y=16'b0000_0100_0000_0000;

		4'b1011:y=16'b0000_1000_0000_0000;

		4'b1100:y=16'b0001_0000_0000_0000;

		4'b1101:y=16'b0010_0000_0000_0000;

		4'b1110:y=16'b0100_0000_0000_0000;

		4'b1111:y=16'b1000_0000_0000_0000;

		default y=16'b0000_0000_0000_0000;
	endcase
end
endmodule
